module lab3_combined(s, o, B, s2, en, R, clock, D, sd);
	parameter N = 32;
	input [4:0] s;
   input [4:0] s2;
	input [4:0]sd; 
	output [N-1:0] B, o;
	wire [N-1:0] m;
	input en;
	input R;
	input clock;
	input [31:0] D;
	
	wire [31:0] Q0, Q1, Q2, Q3, Q4, Q5, Q6, Q7, Q8, Q9, Q10, Q11, Q12, Q13, Q14, Q15, Q16, Q17, Q18, Q19, Q20, Q21, Q22, Q23, Q24, Q25, Q26, Q27, Q28, Q29, Q30, Q31;
	
	lab3_mux instA(o,Q0, Q1, Q2, Q3, Q4, Q5, Q6, Q7, Q8, Q9, Q10, Q11, Q12, Q13, Q14, Q15, Q16, Q17, Q18, Q19, Q20, Q21, Q22, Q23, Q24, Q25, Q26, Q27, Q28, Q29, Q30, Q31, s); 
	lab3_mux instB(B,Q0, Q1, Q2, Q3, Q4, Q5, Q6, Q7, Q8, Q9, Q10, Q11, Q12, Q13, Q14, Q15, Q16, Q17, Q18, Q19, Q20, Q21, Q22, Q23, Q24, Q25, Q26, Q27, Q28, Q29, Q30, Q31, s2); 
	lab3_decoder instX(sd,m, en);
	lab3_register inst0(m[0], Q0, D, R, clock); 
	lab3_register inst1(m[1], Q1, D, R, clock);
	lab3_register inst2(m[2], Q2, D, R, clock);
	lab3_register inst3(m[3], Q3, D, R, clock);
	lab3_register inst4(m[4], Q4, D, R, clock);
	lab3_register inst5(m[5], Q5, D, R, clock);
	lab3_register inst6(m[6], Q6, D, R, clock);
	lab3_register inst7(m[7], Q7, D, R, clock);
	lab3_register inst8(m[8], Q8, D, R, clock);
	lab3_register inst9(m[9], Q9, D, R, clock);
	lab3_register inst10(m[10], Q10, D, R, clock);
	lab3_register inst11(m[11], Q11, D, R, clock);
	lab3_register inst12(m[12], Q12, D, R, clock);
	lab3_register inst13(m[13], Q13, D, R, clock);
	lab3_register inst14(m[14], Q14, D, R, clock);
	lab3_register inst15(m[15], Q15, D, R, clock);
	lab3_register inst16(m[16], Q16, D, R, clock);
	lab3_register inst17(m[17], Q17, D, R, clock);
	lab3_register inst18(m[18], Q18, D, R, clock);
	lab3_register inst19(m[19], Q19, D, R, clock);
	lab3_register inst20(m[20], Q20, D, R, clock);
	lab3_register inst21(m[21], Q21, D, R, clock);
	lab3_register inst22(m[22], Q22, D, R, clock);
	lab3_register inst23(m[23], Q23, D, R, clock);
	lab3_register inst24(m[24], Q24, D, R, clock);
	lab3_register inst25(m[25], Q25, D, R, clock);
	lab3_register inst26(m[26], Q26, D, R, clock);
	lab3_register inst27(m[27], Q27, D, R, clock);
	lab3_register inst28(m[28], Q28, D, R, clock);
	lab3_register inst29(m[29], Q29, D, R, clock);
	lab3_register inst30(m[30], Q30, D, R, clock);
	lab3_register inst31(m[31], Q31, D, R, clock);
endmodule