module lab7_ADD4(in, out4);
	input [7:0] in;
	output [7:0] out4;
	
	assign out4= in + 8'd4;
endmodule
