//decoder
module lab3_decoder(s,m, en); 
	output reg [31:0]m; 
	input [4:0]s; 
	input en;
	
	always @(s or en)   
	begin 
		if (en == 1'b1) 
		case (s) 
			5'b00000: m = 1;
			5'b00001: m = 2;
			5'b00010: m = 4;
			5'b00011: m = 8;
			5'b00100: m = 16;
			5'b00101: m = 32;
			5'b00110: m = 64;
			5'b00111: m = 128;
			5'b01000: m = 256;
			5'b01001: m = 512;
			5'b01010: m = 1024;
			5'b01011: m = 2048;
			5'b01100: m = 4096;
			5'b01101: m = 8192;
			5'b01110: m = 16384;
			5'b01111: m = 32768;
			5'b10000: m = 65536;
			5'b10001: m = 131072;
			5'b10010: m = 262144;
			5'b10011: m = 524288;
			5'b10100: m = 1048576;
			5'b10101: m = 2097152;
			5'b10110: m = 4194304;
			5'b10111: m = 8388608;
			5'b11000: m = 16777216;
			5'b11001: m = 33554432;
			5'b11010: m = 67108864;
			5'b11011: m = 134217728;
			5'b11100: m = 268435456;
			5'b11101: m = 536870912;
			5'b11110: m = 1073741824;
			5'b11111: m = 2147483648;
			default: m = 1'bx; 
		endcase 
		if (en == 0) m = 1'b1; 
	end 
endmodule

